export LANGUAGE="sv_SE.UTF-8"
export LANG="sv_SE.UTF-8"
export LC_ALL="sv_SE.UTF-8"
